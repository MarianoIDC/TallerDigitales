module Suma (A, B, RES, N, Z, C, V);

//Hace cosas de suma
    
endmodule