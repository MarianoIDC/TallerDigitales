module CE();



endmodule 