module OR_Gate ();
    
endmodule