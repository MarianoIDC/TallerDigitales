module Resta ();
    //Hace cosas de Resta
endmodule