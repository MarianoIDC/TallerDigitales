module Modulo ();
    
endmodule