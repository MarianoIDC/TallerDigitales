module Mux #(parameter P=4)();

//Hace cosas de Mux
    
endmodule