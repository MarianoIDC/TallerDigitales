module Multi ();
    //Hace cosas de Multi
    
endmodule