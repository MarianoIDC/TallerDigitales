module RAM_tb();

logic address,
	clock,
	data,
	wren,
	q;


endmodule
