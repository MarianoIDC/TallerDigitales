module Division ();
    // Hace cosas de division 
endmodule