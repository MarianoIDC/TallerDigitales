module CU ();

endmodule
