module sr ();
    
endmodule