module AND_Gate ();
    
endmodule