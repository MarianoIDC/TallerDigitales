module Sumador (input logic [31:0] A, 
					 input logic B,
					 output logic Sum);
					 
		assign Sum = A + B;
		
endmodule 