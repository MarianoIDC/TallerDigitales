module sl ();
    
endmodule