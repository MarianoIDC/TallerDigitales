module XOR_Gate ();
    
endmodule